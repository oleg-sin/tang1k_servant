module toplevel();
endmodule